/* 
* fc_top.v
*/

`timescale 1ns / 1ps

module fc_top 
  #(
    parameter integer C_S00_AXIS_TDATA_WIDTH = 32
  )
  (
    input wire CLK,
    input wire RESETN,

    // AXIS protocol
    output wire S_AXIS_TREADY,
    input wire [C_S00_AXIS_TDATA_WIDTH-1 : 0] S_AXIS_TDATA,
    input wire [(C_S00_AXIS_TDATA_WIDTH/8)-1 : 0] S_AXIS_TKEEP, 
    input wire S_AXIS_TUSER, 
    input wire S_AXIS_TLAST, 
    input wire S_AXIS_TVALID, 

    input wire M_AXIS_TREADY, 
    output wire M_AXIS_TUSER, 
    output wire [C_S00_AXIS_TDATA_WIDTH-1 : 0] M_AXIS_TDATA, 
    output wire [(C_S00_AXIS_TDATA_WIDTH/8)-1 : 0] M_AXIS_TKEEP, 
    output wire M_AXIS_TLAST, 
    output wire M_AXIS_TVALID, 

    // APB protocol
    input wire [31:0] PADDR, 
    input wire PENABLE, 
    input wire PSEL, 
    input wire PWRITE, 
    input wire [31:0] PWDATA, 
    output wire [31:0] PRDATA, 
    output wire PREADY, 
    output wire PSLVERR
  );
  
  // For FC control path
  wire fc_start;
  wire fc_done;
  wire [31:0] clk_counter;
  wire [31:0] max_index;
  assign PREADY = 1'b1;
  assign PSLVERR = 1'b0;

  //////////////////////////////////////////////////////////////////////////
  // [NEW] Wires for Inter-module connection (Command, Status, Config)
  //////////////////////////////////////////////////////////////////////////
  wire [2:0] fc_cmd;           // APB -> Module: Current Command
  wire F_writedone;            // Module -> APB: Status Flag
  wire B_writedone;            // Module -> APB: Status Flag
  wire cal_done;               // Module -> APB: Status Flag
  
  // [NEW] Wires for Variable Size Configuration
  wire [31:0] num_input_words; // APB -> Module: Input Size (FC1/2/3)
  wire [31:0] num_output_words;// APB -> Module: Output Size (FC1/2/3)
  //////////////////////////////////////////////////////////////////////////
  
  clk_counter_fc u_clk_counter(
    .clk   (CLK),
    .rstn  (RESETN),
    .start (fc_start),
    .done  (fc_done),

    .clk_counter (clk_counter)
  );
  
  fc_apb u_fc_apb(
    .PCLK    (CLK),
    .PRESETB (RESETN),
    .PADDR   ({16'd0,PADDR[15:0]}),
    .PSEL    (PSEL),
    .PENABLE (PENABLE),
    .PWRITE  (PWRITE),
    .PWDATA  (PWDATA),
    .PRDATA  (PRDATA),

    .fc_start    (fc_start),
    .fc_done     (fc_done),
    .clk_counter (clk_counter),

    //////////////////////////////////////////////////////////////////////////
    // TODO : Add ports as you need
    //////////////////////////////////////////////////////////////////////////

    .COMMAND          (fc_cmd),           // Output to fc_module
    .F_writedone      (F_writedone),      // Input from fc_module
    .B_writedone      (B_writedone),      // Input from fc_module
    .cal_done         (cal_done),         // Input from fc_module
    .max_index        (max_index),       // Input from fc_module
    
    .num_input_words  (num_input_words),  // Output to fc_module (Register Value)
    .num_output_words (num_output_words)  // Output to fc_module (Register Value)
  );
  
  fc_module u_fc_module(
    .clk  (CLK),
    .rstn (RESETN),

    .S_AXIS_TREADY (S_AXIS_TREADY),
    .S_AXIS_TDATA  (S_AXIS_TDATA),
    .S_AXIS_TKEEP  (S_AXIS_TKEEP),
    .S_AXIS_TUSER  (S_AXIS_TUSER),
    .S_AXIS_TLAST  (S_AXIS_TLAST),
    .S_AXIS_TVALID (S_AXIS_TVALID),

    .M_AXIS_TREADY (M_AXIS_TREADY),
    .M_AXIS_TUSER  (M_AXIS_TUSER),
    .M_AXIS_TDATA  (M_AXIS_TDATA),
    .M_AXIS_TKEEP  (M_AXIS_TKEEP),
    .M_AXIS_TLAST  (M_AXIS_TLAST),
    .M_AXIS_TVALID (M_AXIS_TVALID),

    .fc_start      (fc_start),
    .fc_done       (fc_done),
    //////////////////////////////////////////////////////////////////////////
    // TODO : Add ports as you need
    //////////////////////////////////////////////////////////////////////////
    .COMMAND          (fc_cmd),           // Input Command
    .F_writedone      (F_writedone),      // Output Status
    .B_writedone      (B_writedone),      // Output Status
    .cal_done         (cal_done),         // Output Status
    .max_index        (max_index),        // Output Max Index
    
    .num_input_words  (num_input_words),  // Input Config (Size)
    .num_output_words (num_output_words)  // Input Config (Size)
  );
  
endmodule
